library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity OPERATIONAL_CONTROL_INSTRUCTION_DECODE is
    Port ( R: in STD_LOGIC;
           INSTRUCTION : in STD_LOGIC_VECTOR (15 downto 0);
           CLK : in STD_LOGIC;
           MS : out STD_LOGIC;
           WRITE_REGISTERS : out STD_LOGIC;
           W_ADDRESS : out STD_LOGIC_VECTOR (3 downto 0);
           R_ADDRESS0 : out STD_LOGIC_VECTOR (3 downto 0);
           R_ADDRESS1 : out STD_LOGIC_VECTOR (3 downto 0);
           K : out STD_LOGIC_VECTOR (7 downto 0);
           SR : out STD_LOGIC;
           CT : out STD_LOGIC_VECTOR (3 downto 0);
           KLOAD : out STD_LOGIC;
           INTERNAL_RESET : out STD_LOGIC;
           COND : out STD_LOGIC;
           C : out STD_LOGIC_VECTOR (1 downto 0);
           JUMP : out STD_LOGIC;
           CALL : out STD_LOGIC;
           RET : out STD_LOGIC;
           PORT_CONTROL_ENABLE : out STD_LOGIC;
           PORT_CONTROL_WRITE : out STD_LOGIC);
end OPERATIONAL_CONTROL_INSTRUCTION_DECODE;

architecture OPCONTROLINSTRDECOD of OPERATIONAL_CONTROL_INSTRUCTION_DECODE is

component D_FLIP_FLOP_SYNC_S is
    Port ( D : in STD_LOGIC;
           CLK : in STD_LOGIC;
           S : in STD_LOGIC;
           Q : out STD_LOGIC);
end component;

component DECODER is
    Port ( I : in STD_LOGIC_VECTOR (3 downto 0);
           T : out STD_LOGIC_VECTOR (15 downto 0));
end component;

signal QAUX : STD_LOGIC;
signal TFFQ : STD_LOGIC;
signal INT_R : STD_LOGIC;
signal CTR_CLK : STD_LOGIC := '0';
signal DECODER_OUTPUT : STD_LOGIC_VECTOR (15 downto 0);
signal ALU_OPERATION : STD_LOGIC;
signal ALU_OPERATION_SPECIAL : STD_LOGIC;
signal FLOW_CONTROL_OPERATION : STD_LOGIC;
signal CALL_IN : STD_LOGIC;
signal RET_IN : STD_LOGIC;

begin

FDS0: D_FLIP_FLOP_SYNC_S port map('0', CLK, R, QAUX);
FDS1: D_FLIP_FLOP_SYNC_S port map(QAUX, CLK, R, INT_R);
INTERNAL_RESET <= INT_R;

DCD: DECODER port map(INSTRUCTION(15 downto 12), DECODER_OUTPUT);
ALU_OPERATION_SPECIAL <= DECODER_OUTPUT(13) or DECODER_OUTPUT(12);
ALU_OPERATION <= DECODER_OUTPUT(0) or DECODER_OUTPUT(1) or DECODER_OUTPUT(2) or DECODER_OUTPUT(3) or DECODER_OUTPUT(4) or DECODER_OUTPUT(5) or DECODER_OUTPUT(6) or DECODER_OUTPUT(7) or ALU_OPERATION_SPECIAL;
KLOAD <= (not ALU_OPERATION_SPECIAL and ALU_OPERATION) or DECODER_OUTPUT(14) or DECODER_OUTPUT(10);
WRITE_REGISTERS <= ALU_OPERATION or DECODER_OUTPUT(10) or DECODER_OUTPUT(11);
with ALU_OPERATION_SPECIAL select CT <=
    INSTRUCTION(15 downto 12) when '0',
    INSTRUCTION(3 downto 0) when '1',
    "0000" when others;
SR <= DECODER_OUTPUT(13);
MS <= DECODER_OUTPUT(10) or DECODER_OUTPUT(11);
W_ADDRESS <= INSTRUCTION(11 downto 8);
R_ADDRESS0 <= INSTRUCTION(11 downto 8);
R_ADDRESS1 <= INSTRUCTION(7 downto 4);

FLOW_CONTROL_OPERATION <= DECODER_OUTPUT(9) or DECODER_OUTPUT(8);
COND <= INSTRUCTION(12);
C <= INSTRUCTION(11 downto 10);
JUMP <= (not INSTRUCTION(9)) and INSTRUCTION(8) and FLOW_CONTROL_OPERATION;
CALL <= INSTRUCTION(9) and INSTRUCTION(8) and FLOW_CONTROL_OPERATION;
RET <= (not INSTRUCTION(9)) and (not INSTRUCTION(8)) and INSTRUCTION(7) and (not INSTRUCTION(6))
    and (not INSTRUCTION(5)) and (not INSTRUCTION(4)) and (not INSTRUCTION(3)) and (not INSTRUCTION(3)) 
    and (not INSTRUCTION(2)) and (not INSTRUCTION(1)) and (not INSTRUCTION(0)) and FLOW_CONTROL_OPERATION;
K <= INSTRUCTION(7 downto 0);
PORT_CONTROL_ENABLE <= DECODER_OUTPUT(14) or DECODER_OUTPUT(15) or DECODER_OUTPUT(10) or DECODER_OUTPUT(11);
PORT_CONTROL_WRITE <= DECODER_OUTPUT(14) or DECODER_OUTPUT(15);
end OPCONTROLINSTRDECOD;
